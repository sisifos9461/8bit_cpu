`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date: 2023/05/24 11:18:14
// Design Name: 
// Module Name: store_uni
// Project Name: 
// Target Devices: 
// Tool Versions: 
// Description: 
// 
// Dependencies: 
// 
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
// 
//////////////////////////////////////////////////////////////////////////////////

module store_unit(
    input lm,
    input clk,
    input epr,
    inout [7:0]w
    );
wire [15:0]addr;
mar mar(w[3:0],lm,clk,addr);
prom prom(clk,addr,w,epr);
 
endmodule



module mar(
    input [3:0]win,   //[3:0]w
    input lm,
    input clk,
    output [15:0]out    //prom���
    );
//����
reg [15:0] res;
reg [3:0]in;
always @ (*)
  if(lm) begin
      in = win;
      case(in)
        4'b0000: res = 16'b0000000000000001;
        4'b0001: res = 16'b0000000000000010;
        4'b0010: res = 16'b0000000000000100;
        4'b0011: res = 16'b0000000000001000;
        4'b0100: res = 16'b0000000000010000;
        4'b0101: res = 16'b0000000000100000;
        4'b0110: res = 16'b0000000001000000;
        4'b0111: res = 16'b0000000010000000;
        4'b1000: res = 16'b0000000100000000;
        4'b1001: res = 16'b0000001000000000;
        4'b1010: res = 16'b0000010000000000;
        4'b1011: res = 16'b0000100000000000;
        4'b1100: res = 16'b0001000000000000;
        4'b1101: res = 16'b0010000000000000;
        4'b1110: res = 16'b0100000000000000;
        4'b1111: res = 16'b1000000000000000;
    endcase/*
      res[0] = (in == 4'b0000) ? 1'b1 : 1'b0; // ������Ϊ 0000 ʱ������� 0 λΪ�ߵ�ƽ������λΪ�͵�ƽ
      res[1] = (in == 4'b0001) ? 1'b1 : 1'b0; // ������Ϊ 0001 ʱ������� 1 λΪ�ߵ�ƽ������λΪ�͵�ƽ
      res[2] = (in == 4'b0010) ? 1'b1 : 1'b0; // ������Ϊ 0010 ʱ������� 2 λΪ�ߵ�ƽ������λΪ�͵�ƽ
      res[3] = (in == 4'b0011) ? 1'b1 : 1'b0; // ������Ϊ 0011 ʱ������� 3 λΪ�ߵ�ƽ������λΪ�͵�ƽ
      res[4] = (in == 4'b0100) ? 1'b1 : 1'b0; // ������Ϊ 0100 ʱ������� 4 λΪ�ߵ�ƽ������λΪ�͵�ƽ
      res[5] = (in == 4'b0101) ? 1'b1 : 1'b0; // ������Ϊ 0101 ʱ������� 5 λΪ�ߵ�ƽ������λΪ�͵�ƽ
      res[6] = (in == 4'b0110) ? 1'b1 : 1'b0; // ������Ϊ 0110 ʱ������� 6 λΪ�ߵ�ƽ������λΪ�͵�ƽ
      res[7] = (in == 4'b0111) ? 1'b1 : 1'b0; // ������Ϊ 0111 ʱ������� 7 λΪ�ߵ�ƽ������λΪ�͵�ƽ
      res[8] = (in == 4'b1000) ? 1'b1 : 1'b0; // ������Ϊ 1000 ʱ������� 8 λΪ�ߵ�ƽ������λΪ�͵�ƽ
      res[9] = (in == 4'b1001) ? 1'b1 : 1'b0; // ������Ϊ 1001 ʱ������� 9 λΪ�ߵ�ƽ������λΪ�͵�ƽ
      res[10] = (in == 4'b1010) ? 1'b1 : 1'b0; // ������Ϊ 1010 ʱ������� 10 λΪ�ߵ�ƽ������λΪ�͵�ƽ
      res[11] = (in == 4'b1011) ? 1'b1 : 1'b0; // ������Ϊ 1011 ʱ������� 11 λΪ�ߵ�ƽ������λΪ�͵�ƽ
      res[12] = (in == 4'b1100) ? 1'b1 : 1'b0; // ������Ϊ 1100 ʱ������� 12 λΪ�ߵ�ƽ������λΪ�͵�ƽ
      res[13] = (in == 4'b1101) ? 1'b1 : 1'b0; // ������Ϊ 1101 ʱ������� 13 λΪ�ߵ�ƽ������λΪ�͵�ƽ
      res[14] = (in == 4'b1110) ? 1'b1 : 1'b0; // ������Ϊ 1110 ʱ������� 14 λΪ�ߵ�ƽ������λΪ�͵�ƽ
      res[15] = (in == 4'b1111) ? 1'b1 : 1'b0; // ������Ϊ 1111 ʱ������� 15 λΪ�ߵ�ƽ������λΪ�͵�ƽ
  */end  
  else begin
     in = 4'hz;
     res = 16'hzzzz;
  end

assign out = res;
endmodule

module prom (
    input clk,         // ʱ���ź�
    input [15:0]addr,  // ��ַ�źţ�16 λ��������
    output[7:0]inst,  // �洢����ָ��������8 λ��������  ��������w
    input epr
);

reg [7:0]reinst;
//reg [7:0] mem [0:255]; // ����һ�� 256 �� 8 λԪ�صĴ洢��
reg [7:0]mem[0:15];
integer j;
integer i;

always @(posedge clk)
   case(addr)
        16'b0000000000000001: reinst =8'b00001111;  //0
        16'b0000000000000010: reinst= 8'b11100000;  //e
        16'b0000000000000100: reinst= 8'b00001111;   //0
        16'b0000000000001000: reinst= 8'b00111110;   //3
        16'b0000000000010000: reinst= 8'b11100000;  //e
        16'b0000000000100000: reinst= 8'b01101101;  //6
        16'b0000000001000000: reinst= 8'b01110011; //7
        16'b0000000010000000: reinst= 8'b11110000;   //f
        16'b0000000100000000: reinst= 8'b00000000;
        16'b0000001000000000: reinst= 8'b00000000;
        16'b0000010000000000: reinst= 8'b00000000;
        16'b0000100000000000: reinst= 8'b00000000;
        16'b0001000000000000: reinst= 8'b00000000;
        16'b0010000000000000: reinst= 8'b00010000;  //16
        16'b0100000000000000: reinst= 8'b00000010; //2
        16'b1000000000000000: reinst= 8'b00000001; //1
    endcase     
assign inst = (epr)?reinst: 8'hzz;
        
        
/*
initial begin
    mem[0] = 8'b00001111;  // MOV ��,(RF)
    mem[1] = 8'b00111110;  // ADD A, (RE)
    mem[2] = 8'b1110xxxx;  // OUT(n),A
    mem[3] = 8'b1111xxxx;  //CPU��ͣ
    for (j = 4; j <14; j = j + 1) begin
      mem[i] = 8'b00000000;
    end
    mem[14] = 8'b00100000;   //32
    mem[15] = 8'b01000000;   //64
    
      
    
end

always @* 
    for(i=0;i<16;i=i+1)begin
         //$display($realtime,"%b,%b,%b,%b,%b",i,reinst,addr[i],addr,inst);
        if(addr[i])begin
            reinst = mem[i]; // ���洢���ж�Ӧ��ַ��ָ�����
        end
    end


assign inst = (epr)?reinst: 8'hzz;
*/
endmodule

